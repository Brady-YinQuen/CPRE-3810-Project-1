library IEEE;
use IEEE.std_logic_1164.all;

entity n_reg_tb is
    generic(gCLK_HPER   : time := 50 ns;
    		N : integer := 32);
end n_reg_tb;

architecture behavior of n_reg_tb is

    constant cCLK_PER  : time := gCLK_HPER * 2;

    component N_Reg is port(
        i_CLK        : in std_logic;  
        i_RST        : in std_logic;
        i_WE         : in std_logic;
        i_D          : in std_logic_vector(N-1 downto 0);
        o_Q          : out std_logic_vector(N-1 downto 0)
        );
    end component;

    signal s_CLK, s_RST, s_WE : std_logic;
    signal s_D, s_Q : std_logic_vector(N-1 downto 0);

begin
    REG_Nbit : N_Reg 
    port map(
        i_CLK   => s_CLK,
        i_RST   => s_RST,
        i_WE    => s_WE,
        i_D     => s_D,
        o_Q     => s_Q
    );

    stimulus_process: process
    begin
        s_CLK <= '0';
        wait for gCLK_HPER;
        s_CLK <= '1';
        wait for gCLK_HPER;
    end process;

    tb_process: process
    begin
        -- Reset the FF
        s_RST <= '1';
        s_WE  <= '0';
        s_D   <= x"00000000";
        wait for cCLK_PER;
    
        -- Store 'FFFFFFFF'
        s_RST <= '0';
        s_WE  <= '1';
        s_D   <= x"FFFFFFFF";
        wait for cCLK_PER;  
    
        -- Keep 'FFFFFFFFF'
        s_RST <= '0';
        s_WE  <= '0';
        s_D   <= x"00000000";
        wait for cCLK_PER;  
    
        -- Store '0'    
        s_RST <= '0';
        s_WE  <= '1';
        s_D   <= x"00000000";
        wait for cCLK_PER;  
    
        -- Keep '0'
        s_RST <= '0';
        s_WE  <= '0';
        s_D   <= x"FFFFFFFF";
        wait for cCLK_PER;  

    end process;



end behavior ; 