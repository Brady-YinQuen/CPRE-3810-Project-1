library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all; -- For arithmetic on std_logic_vector

entity N_decoder is
    generic(N : integer := 5);  -- N is 5 for a 5-bit decoder
    port(
        i_sel : in std_logic_vector(N-1 downto 0);
        o_O   : out std_logic_vector(2**N-1 downto 0)  -- Output of size 32-bits
    );
end N_decoder;

architecture dataflow of N_decoder is
begin
with i_sel select

o_O  <= x"00000001" when "00000",
	x"00000002" when "00001",  -- bit 1 set
       x"00000004" when "00010",  -- bit 2 set
       x"00000008" when "00011",  -- bit 3 set
       x"00000010" when "00100",  -- bit 4 set
       x"00000020" when "00101",  -- bit 5 set
       x"00000040" when "00110",  -- bit 6 set
       x"00000080" when "00111",  -- bit 7 set
       x"00000100" when "01000",  -- bit 8 set
       x"00000200" when "01001",  -- bit 9 set
       x"00000400" when "01010",  -- bit 10 set
       x"00000800" when "01011",  -- bit 11 set
       x"00001000" when "01100",  -- bit 12 set
       x"00002000" when "01101",  -- bit 13 set
       x"00004000" when "01110",  -- bit 14 set
       x"00008000" when "01111",  -- bit 15 set
       x"00010000" when "10000",  -- bit 16 set
       x"00020000" when "10001",  -- bit 17 set
       x"00040000" when "10010",  -- bit 18 set
       x"00080000" when "10011",  -- bit 19 set
       x"00100000" when "10100",  -- bit 20 set
       x"00200000" when "10101",  -- bit 21 set
       x"00400000" when "10110",  -- bit 22 set
       x"00800000" when "10111",  -- bit 23 set
       x"01000000" when "11000",  -- bit 24 set
       x"02000000" when "11001",  -- bit 25 set
       x"04000000" when "11010",  -- bit 26 set
       x"08000000" when "11011",  -- bit 27 set
       x"10000000" when "11100",  -- bit 28 set
       x"20000000" when "11101",  -- bit 29 set
       x"40000000" when "11110",  -- bit 30 set
       x"80000000" when "11111",   -- bit 31 set
	x"00000000" when others;

end dataflow;