library IEEE;
use IEEE.std_logic_1164.all;
use work.my_package.all;

entity MIP_REG_tb is
    generic(gCLK_HPER   : time := 50 ns);
end entity MIP_REG_tb;

architecture behavior of MIP_REG_tb is
    constant cCLK_PER  : time := gCLK_HPER * 2;
    component MIP_REG is
        port(
            i_rs : in std_logic_vector(4 downto 0);
            i_rt : in std_logic_vector(4 downto 0);
            i_rd : in std_logic_vector(4 downto 0);
            i_d  : in std_logic_vector(31 downto 0);
            i_reset : in std_logic;  
            i_clock : in std_logic;  
            i_we    : in std_logic;
            o_D1    : out std_logic_vector(31 downto 0);
            o_D2    : out std_logic_vector(31 downto 0)
        );
    end component MIP_REG;

    signal s_rs :  std_logic_vector(4 downto 0);
    signal s_rt :  std_logic_vector(4 downto 0);
    signal s_rd :  std_logic_vector(4 downto 0);
    signal s_d  :  std_logic_vector(31 downto 0);
    signal s_reset :  std_logic;  
    signal s_clock :  std_logic;  
    signal s_we    :  std_logic;
    signal s_D1    :  std_logic_vector(31 downto 0);
    signal s_D2    :  std_logic_vector(31 downto 0);

    begin 
        g_Mip : MIP_REG
        port map(
            i_rs => s_rs,
            i_rt => s_rt,
            i_rd => s_rd,
            i_d  => s_d,
            i_reset => s_reset,
            i_clock => s_clock,  
            i_we    => s_we,
            o_D1    => s_D1,
            o_D2    => s_D2
        );

        stimulus_process: process
        begin
            s_clock <= '0';
            wait for gCLK_HPER;
            s_clock <= '1';
            wait for gCLK_HPER;
        end process;

        simulation: process
        begin 
        s_reset <= '1';
        s_we <= '1';
        s_rs <= "00000";
        s_rt <= "00000";
        s_rd <= "00000";
        s_d  <= x"00000000";
        wait for cCLK_PER;


        s_reset <= '0';
        s_we <= '1' ;
        s_rs <= "00000";
        s_rt <= "00001";
        s_rd <= "00000";
        s_d  <= x"FFFFFFFF";
        wait for cCLK_PER;

 	s_reset <= '0';
        s_we <= '1' ;
        s_rs <= "00000";
        s_rt <= "00001";
        s_rd <= "00001";
        s_d  <= x"0BEFACED";
        wait for cCLK_PER;

    end process;





end architecture behavior;