library IEEE;
use IEEE.std_logic_1164.all;
use work.my_package.all;

entity MySecondMIPSDatapath_tb is
    generic(gCLK_HPER   : time := 10 ns);
end entity MySecondMIPSDatapath_tb;

architecture behavior of MySecondMIPSDatapath_tb  is
    constant cCLK_PER  : time := gCLK_HPER * 2;
    component MySecondMIPSDatapath is
        port (
            i_rs : in std_logic_vector(4 downto 0);
            i_rt : in std_logic_vector(4 downto 0);
            i_rd : in std_logic_vector(4 downto 0);
            i_reset : in std_logic;  
            i_clock : in std_logic;  
            i_we    : in std_logic; 
            i_addsub_en : in std_logic;   -- this is to select add or sub 
            i_imm: in  std_logic_vector(15 downto 0);
            i_ALUSrc : in std_logic;
            i_sw_en : in std_logic;
            i_sign_ext : in std_logic;
            i_memToReg_en : in std_logic;
            o_OF : out std_logic;
            o_ALU_debug: out std_logic_vector(31 downto 0)
        );
        end component MySecondMIPSDatapath;

        signal s_rs :  std_logic_vector(4 downto 0);
        signal s_rt :  std_logic_vector(4 downto 0);
        signal s_rd :  std_logic_vector(4 downto 0);
        signal s_reset  :  std_logic;  
        signal s_clock  :  std_logic;  
        signal s_we     :  std_logic;
        signal s_addsub_en :  std_logic; 
        signal s_imm    :  std_logic_vector(15 downto 0);
        signal s_ALUSrc :  std_logic;
        signal s_sw_en  :  std_logic;
        signal s_sign_ext : std_logic;
        signal s_memToReg_en : std_logic;
        signal s_OF     :  std_logic;
	    signal s_ALU_debug:  std_logic_vector(31 downto 0);

        begin
            g_mip_alu: MySecondMIPSDatapath
            port Map(
                i_rs    => s_rs,
                i_rt    => s_rt,
                i_rd    => s_rd,
                i_reset => s_reset,
                i_clock => s_clock,  
                i_we    => s_we,
                i_addsub_en     => s_addsub_en,
                i_imm           => s_imm,
                i_ALUSrc        => s_ALUSrc,  
                i_sw_en         => s_sw_en,
                i_sign_ext      => s_sign_ext, 
                i_memToReg_en   => s_memToReg_en, 
                o_OF            => s_OF,
                o_ALU_debug     => s_ALU_debug
            );


            stimulus_process: process
            begin
                s_clock <= '0';
                wait for gCLK_HPER;
                s_clock <= '1';
                wait for gCLK_HPER;
            end process;

            simulation: process
            begin

                s_reset <= '1';
                wait for cCLK_PER;
                s_reset <= '0';
                wait for cCLK_PER;

	--	s_rs <= "00000";
    --            s_rt <= "00000";
    --            s_rd <= "00001";
     --           s_we    <= '1';
  --              s_addsub_en     <= '0';
     --           s_imm   <=  x"0005";
   --             s_ALUSrc  <= '1';  
     --           s_sw_en <= '0';
   --             s_sign_ext <= '0';
  --              s_memToReg_en <= '0';
  --              wait for cCLK_PER;
--
	--	s_rs <= "00000";
  --              s_rt <= "00001";
   --             s_rd <= "00001";
  --              s_we    <= '0';
  --              s_addsub_en     <= '0';
 --               s_imm   <=  x"0000";
  --              s_ALUSrc  <= '1';  
  --              s_sw_en <= '1';
  --              s_sign_ext <= '0';
    --            s_memToReg_en <= '0';
  --              wait for cCLK_PER;

	--	s_rs <= "00000";
 --               s_rt <= "00001";
--                s_rd <= "00010";
 --               s_we    <= '1';
--                s_addsub_en     <= '0';
 --               s_imm   <=  x"0000";
 --               s_ALUSrc  <= '1';  
 --               s_sw_en <= '0';
  --              s_sign_ext <= '0';
 --               s_memToReg_en <= '1';
 --               wait for cCLK_PER;



                -- case 1
                s_rs <= "00000";
                s_rt <= "00000";
                s_rd <= "11001";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0000";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

                -- case 2
                s_rs <= "00000";
                s_rt <= "00000";
                s_rd <= "11010";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0100";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 3
                s_rs <= "11001";
                s_rt <= "00000";
                s_rd <= "00001";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0000";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '1';
                wait for cCLK_PER;
		
		-- case 4
                s_rs <= "11001";
                s_rt <= "00000";
                s_rd <= "00010";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '1';
                wait for cCLK_PER;

		-- case 5 expected 6 
		s_rs <= "00001";
                s_rt <= "00010";
                s_rd <= "00001";
                s_we    <= '1';
                s_addsub_en    <= '0';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '0';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		
		-- case 6 storing 6 to 256mem
		s_rs <= "11010";
                s_rt <= "00001";
                s_rd <= "00001";
                s_we    <= '0';
                s_addsub_en     <= '0';
                s_imm   <=  x"0000";
                s_ALUSrc  <= '1';  
                s_sw_en <= '1';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 7
                s_rs <= "11001";
                s_rt <= "00000";
                s_rd <= "00010";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0008";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '1';
                wait for cCLK_PER;

		-- case 8 expected F
		s_rs <= "00001";
                s_rt <= "00010";
                s_rd <= "00001";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '0';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 9 storing F to 256 + 4 mem
		s_rs <= "11010";
                s_rt <= "00001";
                s_rd <= "00001";
                s_we    <= '0';
                s_addsub_en     <= '0';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '1';  
                s_sw_en <= '1';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 10 
                s_rs <= "11001";
                s_rt <= "00000";
                s_rd <= "00010";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"000C";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '1';
                wait for cCLK_PER;
		


		-- case 11 expected is 1b
		s_rs <= "00001";
                s_rt <= "00010";
                s_rd <= "00001";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '0';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 12 storing 1B to 256 + 4 mem
		s_rs <= "11010";
                s_rt <= "00001";
                s_rd <= "00001";
                s_we    <= '0';
                s_addsub_en     <= '0';
                s_imm   <=  x"0008";
                s_ALUSrc  <= '1';  
                s_sw_en <= '1';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;


		-- case 13 
                s_rs <= "11001";
                s_rt <= "00000";
                s_rd <= "00010";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0010";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '1';
                wait for cCLK_PER;

		-- case 14 expected is 1d
		s_rs <= "00001";
                s_rt <= "00010";
                s_rd <= "00001";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '0';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 15 storing 1d to 256 + 4 mem
		s_rs <= "11010";
                s_rt <= "00001";
                s_rd <= "00001";
                s_we    <= '0';
                s_addsub_en     <= '0';
                s_imm   <=  x"000C";
                s_ALUSrc  <= '1';  
                s_sw_en <= '1';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 16 
                s_rs <= "11001";
                s_rt <= "00000";
                s_rd <= "00010";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0014";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '1';
                wait for cCLK_PER;

		-- case 17 expected is 23
		s_rs <= "00001";
                s_rt <= "00010";
                s_rd <= "00001";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '0';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 18 storing 23 to 256 + 4 mem
		s_rs <= "11010";
                s_rt <= "00001";
                s_rd <= "00001";
                s_we    <= '0';
                s_addsub_en     <= '0';
                s_imm   <=  x"0010";
                s_ALUSrc  <= '1';  
                s_sw_en <= '1';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 19 
                s_rs <= "11001";
                s_rt <= "00000";
                s_rd <= "00010";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0018";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '1';
                wait for cCLK_PER;

		-- case 20 expected is 2d
		s_rs <= "00001";
                s_rt <= "00010";
                s_rd <= "00001";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '0';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;

		-- case 21 
		s_rs <= "00000";
                s_rt <= "00010";
                s_rd <= "11011";
                s_we    <= '1';
                s_addsub_en     <= '0';
                s_imm   <=  x"0200";
                s_ALUSrc  <= '1';  
                s_sw_en <= '0';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;


		-- case 22 
		s_rs <= "11011";
                s_rt <= "00001";
                s_rd <= "00001";
                s_we    <= '0';
                s_addsub_en     <= '1';
                s_imm   <=  x"0004";
                s_ALUSrc  <= '1';  
                s_sw_en <= '1';
                s_sign_ext <= '0';
                s_memToReg_en <= '0';
                wait for cCLK_PER;


		


                 

            end process;







        end architecture behavior ; 