library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_Shifter is
end tb_Shifter;

architecture behavior of tb_Shifter is

    component Shifter is 
    port(
        i_shiftamount: in std_logic_vector(4 downto 0);
        i_data: in std_logic_vector(31 downto 0);
        i_shiftright: in std_logic;
        i_arithmetic: in std_logic;
        o_data: out std_logic_vector(31 downto 0)
    );
    end component Shifter;


    signal s_shiftamount : std_logic_vector(4 downto 0);
    signal s_data        : std_logic_vector(31 downto 0);
    signal s_shiftright   : std_logic;
    signal s_arithmetic  : std_logic;
    signal s_o_data        : std_logic_vector(31 downto 0);
begin
    -- Instantiate the Shifter
    uut: Shifter
        port map(
            i_shiftamount => s_shiftamount,
            i_data        => s_data,
            i_shiftright   => s_shiftright,
            i_arithmetic  => s_arithmetic,
            o_data        => s_o_data
        );

    -- Test process
    process
    begin
        -- Test case 1: Shift right by FFFFFFF
        s_data <= x"10101010";
        s_shiftamount <= "11111";
        s_shiftright <= '1';
        s_arithmetic <= '0';
        wait for 10 ns;

        -- Test case 2: Logical shift right by 3
        s_data <= x"00000001";
        s_shiftamount <= "00011";
        s_shiftright <= '1';
        s_arithmetic <= '0';
        wait for 10 ns;
   

        -- Test case 3: Arithmetic shift right by 1
        s_data <= x"00000008";
        s_shiftamount <= "00010";
        s_shiftright <= '1';
        s_arithmetic <= '1';
        wait for 10 ns;
  

        wait;
    end process;
end behavior;